module ssss
ssss
endmodule